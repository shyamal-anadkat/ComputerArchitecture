module xor2(a, b, out);
	input a, b; 
	output out; 
	assign Out = a ^ b;
endmodule 
