module cla16 (A, B, Cin, Cout, PG, GG, S);

   input [15:0] A, B;
   input Cin;
   output [15:0] S;
   output Cout, PG, GG;

   wire [15:0] G, P, C; 

endmodule