module ripple_4 (
	input [3:0] A, B,
	output [3:0] SUM );



endmodule
