module xor2(In1, In2, Out);
	input In1, In2; 
	output Out; 
	assign Out = In1^In2; 
endmodule 